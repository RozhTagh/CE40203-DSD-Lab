library verilog;
use verilog.vl_types.all;
entity booth_TB is
end booth_TB;
